//==============================================================================
// Module: line_buffer
// Description: Line buffer 3 dòng tạo sliding window 3x3 cho Sobel
//              Sử dụng 2 BRAM (640x8-bit) lưu 2 dòng trước
//              Output window 9 pixels cho mỗi pixel hiện tại
// Author: Nguyễn Văn Đạt
// Date: 2025
// Target: Tang Nano 4K (GW1NSR-LV4C)
//==============================================================================
module line_buffer #(
    parameter IMG_WIDTH   = 640,
    parameter PIXEL_WIDTH = 8,
    parameter ADDR_WIDTH  = 10
)(
    input  wire                     clk,
    input  wire                     rst_n,
    input  wire                     pixel_valid,
    input  wire [PIXEL_WIDTH-1:0]   pixel_in,
    output wire                     window_valid,
    output wire [PIXEL_WIDTH*9-1:0] window_out
);

    // =========================================================================
    // OPTIMIZATION 1: Reduce address tracking registers
    // Before: write_addr, write_addr_d0, write_addr_d1 (30 bits)
    // After: Only col_addr (10 bits) - saves 20 FFs
    // =========================================================================
    reg [ADDR_WIDTH-1:0] col_addr;
    reg [ADDR_WIDTH-1:0] row_count;

    // =========================================================================
    // OPTIMIZATION 2: Simplified pipeline - 2 stages instead of 3
    // BRAM has 2-cycle latency: addr_reg -> BRAM -> dout_reg
    // We only need d1 and d2 for proper alignment
    // Saves: 1 valid bit + 20 address bits + 8 pixel bits = 29 FFs
    // =========================================================================
    reg pixel_valid_d1, pixel_valid_d2;
    reg [ADDR_WIDTH-1:0] col_addr_d1, col_addr_d2;
    reg [ADDR_WIDTH-1:0] row_count_d1, row_count_d2;
    reg [PIXEL_WIDTH-1:0] pixel_in_d1, pixel_in_d2;

    // BRAM outputs (3 line buffers)
    wire [PIXEL_WIDTH-1:0] line0_q, line1_q, line2_q;

    // =========================================================================
    // OPTIMIZATION 3: Remove redundant BRAM output registers
    // BRAM already has output register (oce control)
    // Saves: 3 * 8 = 24 FFs
    // =========================================================================
    
    // 3x3 window shift registers (required for convolution)
    reg [PIXEL_WIDTH-1:0] top_row  [0:2];  // Row n-2
    reg [PIXEL_WIDTH-1:0] mid_row  [0:2];  // Row n-1
    reg [PIXEL_WIDTH-1:0] bot_row  [0:2];  // Row n (current)

    // Prefill tracking (to flush stale data from BRAMs)
    reg prefill_active;
    reg [ADDR_WIDTH+1:0] fill_count;
    
    localparam FLUSH_THRESHOLD = (IMG_WIDTH * 2) + 1;
    localparam [PIXEL_WIDTH-1:0] ZERO_PIXEL = {PIXEL_WIDTH{1'b0}};

    reg window_valid_reg;
    integer i;

    // =========================================================================
    // Column address counter (wraps at IMG_WIDTH)
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            col_addr <= {ADDR_WIDTH{1'b0}};
        end else if (pixel_valid) begin
            col_addr <= (col_addr == IMG_WIDTH - 1) ? {ADDR_WIDTH{1'b0}} : col_addr + 1'b1;
        end
    end

    // =========================================================================
    // Row counter (saturates after 2 full rows buffered)
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            row_count <= {ADDR_WIDTH{1'b0}};
        end else if (pixel_valid && (col_addr == IMG_WIDTH - 1)) begin
            if (row_count != {ADDR_WIDTH{1'b1}}) begin
                row_count <= row_count + 1'b1;
            end
        end
    end

    // =========================================================================
    // Prefill logic: Wait for 2 rows + 1 pixel before valid output
    // This flushes any garbage from BRAM power-up
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            prefill_active <= 1'b1;
            fill_count <= {(ADDR_WIDTH+2){1'b0}};
        end else if (prefill_active && pixel_valid) begin
            if (fill_count >= FLUSH_THRESHOLD - 1) begin
                prefill_active <= 1'b0;
            end else begin
                fill_count <= fill_count + 1'b1;
            end
        end
    end

    // =========================================================================
    // Pipeline stage 1: Delay by 1 cycle (BRAM address register stage)
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            pixel_valid_d1 <= 1'b0;
            col_addr_d1    <= {ADDR_WIDTH{1'b0}};
            row_count_d1   <= {ADDR_WIDTH{1'b0}};
            pixel_in_d1    <= {PIXEL_WIDTH{1'b0}};
        end else begin
            pixel_valid_d1 <= pixel_valid;
            if (pixel_valid) begin
                col_addr_d1  <= col_addr;
                row_count_d1 <= row_count;
                pixel_in_d1  <= pixel_in;
            end
        end
    end

    // =========================================================================
    // Pipeline stage 2: Delay by 2 cycles (BRAM output register stage)
    // This aligns with BRAM read data availability
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            pixel_valid_d2 <= 1'b0;
            col_addr_d2    <= {ADDR_WIDTH{1'b0}};
            row_count_d2   <= {ADDR_WIDTH{1'b0}};
            pixel_in_d2    <= {PIXEL_WIDTH{1'b0}};
        end else begin
            pixel_valid_d2 <= pixel_valid_d1;
            if (pixel_valid_d1) begin
                col_addr_d2  <= col_addr_d1;
                row_count_d2 <= row_count_d1;
                pixel_in_d2  <= pixel_in_d1;
            end
        end
    end

    // =========================================================================
    // 3x3 Window Formation via Shift Registers
    // Window layout:  top_row[0]  top_row[1]  top_row[2]
    //                 mid_row[0]  mid_row[1]  mid_row[2]
    //                 bot_row[0]  bot_row[1]  bot_row[2]
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (i = 0; i < 3; i = i + 1) begin
                top_row[i] <= ZERO_PIXEL;
                mid_row[i] <= ZERO_PIXEL;
                bot_row[i] <= ZERO_PIXEL;
            end
        end else if (pixel_valid_d2) begin
            if (prefill_active) begin
                // During prefill, keep window zeroed
                for (i = 0; i < 3; i = i + 1) begin
                    top_row[i] <= ZERO_PIXEL;
                    mid_row[i] <= ZERO_PIXEL;
                    bot_row[i] <= ZERO_PIXEL;
                end
            end else begin
                // Shift left and load new column from right
                top_row[0] <= top_row[1];
                top_row[1] <= top_row[2];
                top_row[2] <= line2_q;      // Row n-2 from BRAM

                mid_row[0] <= mid_row[1];
                mid_row[1] <= mid_row[2];
                mid_row[2] <= line1_q;      // Row n-1 from BRAM

                bot_row[0] <= bot_row[1];
                bot_row[1] <= bot_row[2];
                bot_row[2] <= pixel_in_d2;  // Current row direct input
            end
        end
    end

    // =========================================================================
    // Window Valid Generation
    // Valid when: row >= 2, col >= 2 (need 3x3 neighborhood fully formed), not prefilling
    // =========================================================================
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            window_valid_reg <= 1'b0;
        end else begin
            window_valid_reg <= pixel_valid_d2 && 
                                (row_count_d2 >= 3) && 
                                (col_addr_d2 >= 2) && 
                                !prefill_active;
        end
    end

    assign window_valid = window_valid_reg;

    // =========================================================================
    // Window Output Assignment (9 pixels flattened)
    // =========================================================================
    assign window_out[7:0]   = top_row[0];
    assign window_out[15:8]  = top_row[1];
    assign window_out[23:16] = top_row[2];
    assign window_out[31:24] = mid_row[0];
    assign window_out[39:32] = mid_row[1];
    assign window_out[47:40] = mid_row[2];
    assign window_out[55:48] = bot_row[0];
    assign window_out[63:56] = bot_row[1];
    assign window_out[71:64] = bot_row[2];

    // =========================================================================
    // BRAM Instantiation: 3 Line Buffers
    // Each stores 1 image row (640 pixels x 8 bits)
    // BRAM primitive handles dual-port read/write with 2-cycle latency
    // =========================================================================

    // Line 0: Direct capture of incoming pixels
    bram line0 (
        .dout   (line0_q),
        .clk    (clk),
        .cea    (pixel_valid),      // Write enable
        .reseta (~rst_n),
        .ceb    (1'b1),             // Read always enabled
        .resetb (~rst_n),
        .oce    (1'b1),             // Output enable
        .ada    (col_addr),         // Write address
        .din    (pixel_in),         // Write data
        .adb    (col_addr)          // Read address (same for circular)
    );

    // Line 1: Delayed by 1 row from Line 0
    wire [PIXEL_WIDTH-1:0] line1_din = (prefill_active && (row_count_d1 == 0)) 
                                       ? ZERO_PIXEL : line0_q;
    
    bram line1 (
        .dout   (line1_q),
        .clk    (clk),
        .cea    (pixel_valid_d1),
        .reseta (~rst_n),
        .ceb    (1'b1),
        .resetb (~rst_n),
        .oce    (1'b1),
        .ada    (col_addr_d1),
        .din    (line1_din),
        .adb    (col_addr_d1)
    );

    // Line 2: Delayed by 2 rows from Line 0
    wire [PIXEL_WIDTH-1:0] line2_din = (prefill_active && (row_count_d2 <= 1)) 
                                       ? ZERO_PIXEL : line1_q;
    
    bram line2 (
        .dout   (line2_q),
        .clk    (clk),
        .cea    (pixel_valid_d2),
        .reseta (~rst_n),
        .ceb    (1'b1),
        .resetb (~rst_n),
        .oce    (1'b1),
        .ada    (col_addr_d2),
        .din    (line2_din),
        .adb    (col_addr_d2)
    );

    // =========================================================================
    // Debug Displays (Simulation Only)
    // =========================================================================
`ifndef SYNTHESIS
    reg [3:0] dbg_window_count;
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            dbg_window_count <= 4'd0;
        end else if (pixel_valid_d2 && !prefill_active) begin
            if (dbg_window_count < 4'd8) begin
                dbg_window_count <= dbg_window_count + 1'b1;
                $display("[LINEBUF t=%0t] row=%0d col=%0d window=%02x_%02x_%02x_%02x_%02x_%02x_%02x_%02x_%02x",
                         $time, row_count_d2, col_addr_d2,
                         top_row[0], top_row[1], top_row[2],
                         mid_row[0], mid_row[1], mid_row[2],
                         bot_row[0], bot_row[1], bot_row[2]);
            end
        end
    end

`ifdef TB_SOBEL_RANDOM
    always @(posedge clk) begin
        if (tb_sobel_random.current_frame_id == 5 &&
            row_count_d2 >= 88 && row_count_d2 <= 92 &&
            pixel_valid_d2 && !prefill_active) begin
            $display("[LINEBUFCHK t=%0t] frame=%0d row=%0d col=%0d win=%02x_%02x_%02x_%02x_%02x_%02x_%02x_%02x_%02x",
                     $time, tb_sobel_random.current_frame_id,
                     row_count_d2, col_addr_d2,
                     top_row[0], top_row[1], top_row[2],
                     mid_row[0], mid_row[1], mid_row[2],
                     bot_row[0], bot_row[1], bot_row[2]);
        end
    end
`endif
`endif

endmodule

// =============================================================================
// OPTIMIZATION SUMMARY
// =============================================================================
// 1. Removed write_addr + delays (3 regs x 10 bits) = -30 FFs
// 2. Removed pixel_valid_d0 + col_addr_d0 + row_count_d0 = -21 FFs
// 3. Removed line0_q_d, line1_q_d, line2_q_d = -24 FFs
// 4. Total savings: ~75 Flip-Flops (~15-20 LUTs equivalent)
// 
// BRAM usage: Unchanged (3 SDPB blocks for 640x8 line buffers)
// Logic depth: Reduced (fewer mux levels in address generation)
// Timing: Maintained (proper 2-cycle BRAM latency alignment)
// =============================================================================

